
module part2(input logic Clock, Reset_b, input logic[ 7:0] Data, input logic [1:0] Function, input logic [7:0] ALUout);
