module part3(input logic clock, input logic reset, ParallelLoadn, RotateRight, ASRight, Data_IN, Q);


